--Sprites
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.numeric_std.all;


use work.game_board_array.all;
use work.Sprite_set.all;
use work.Sprite_Image.all;
use work.game_board_free.all;
use work.standard_sprite.all;


entity Sprites is
	Port (
			Reset : in std_logic;
			DrawX : in std_logic_vector (9 downto 0);
			DrawY : in std_logic_vector (9 downto 0);
			outFree : in game_board_free_spaces;
			outSprites: in sprite_location;
			scoreIn : in scoreBoard;
			--sprite_img : out img;
			sprite_num_color : out std_logic_vector (29 downto 0);
			sprite_back_color : out std_logic_vector (29 downto 0);
			tile_sprite_out : out img;
			score_sprite_out : out array_16x16);

end Sprites;

architecture Behavioral of Sprites is

	
	--type array_16x16 is array (0 to 15) of std_logic_vector (15 downto 0);
	constant sprite_S : array_16x16 := 
		("0000000000000000", --capital S
		 "0000000000000000",
		 "0000000000000000",
		 "0000111111111000",
		 "0001111111111000",
		 "0001100000000000",
		 "0001100000000000",
		 "0001111111111000",
		 "0000111111111000",
		 "0000000000011000",
		 "0000000000011000",
		 "0001111111111000",
		 "0001111111110000",
		 "0000000000000000",
		 "0000000000000000",
		 "0000000000000000");
	constant sprite_C : array_16x16 := 
		("0000000000000000", --capital C
		"0000000000000000", 
	    "0000000000000000", 
		"0000111111111000", 
		"0001111111111000", 
		"0001100000000000", 
		"0001100000000000", 
		"0001100000000000", 
		"0001100000000000", 
		"0001100000000000", 
		"0001100000000000", 
		"0001111111111000", 
		"0000111111111000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_O : array_16x16 := 
		("0000000000000000", --capital O
		"0000000000000000", 
		"0000000000000000", 
		"0000111111110000", 
		"0001111111111000", 
		"0001100000011000", 
		"0001100000011000", 
		"0001100000011000", 
		"0001100000011000", 
		"0001100000011000", 
		"0001100000011000", 
		"0001111111111000", 
		"0000111111110000", 
		"0000000000000000",
		"0000000000000000", 
		"0000000000000000");
	constant sprite_R : array_16x16 := 
		("0000000000000000", --capital R
		"0000000000000000", 
		"0000000000000000", 
		"0000111111110000", 
		"0001111111111000", 
		"0001100000011000", 
		"0001100000011000", 
		"0001111111111000", 
		"0001111111110000", 
		"0001100111000000", 
		"0001100011100000", 
		"0001100001110000", 
		"0001100000111000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_E : array_16x16 :=
		("0000000000000000", --capital E
		"0000000000000000", 
		"0000000000000000", 
		"0001111111111000", 
		"0001111111111000", 
		"0001100000000000", 
		"0001100000000000", 
		"0001111111111000", 
		"0001111111111000", 
		"0001100000000000", 
		"0001100000000000", 
		"0001111111111000", 
		"0001111111111000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	
	constant sprite_score_0	: array_16x16 :=
		("0000000000000000", --0 used for keeping score
		"0000000000000000", 
		"0000000000000000", 
		"0000111111110000", 
		"0001111111111000", 
		"0001100000111000", 
		"0001100001011000", 
		"0001100010011000", 
		"0001100100011000", 
		"0001101000011000", 
		"0001110000011000", 
		"0001111111111000", 
		"0000111111110000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_score_1	: array_16x16 :=
		("0000000000000000", --1 used for keeping score
		"0000000000000000", 
		"0000000000000000", 
		"0000001111000000", 
		"0000011111000000", 
		"0000111111000000", 
		"0000000111000000", 
		"0000000111000000", 
		"0000000111000000", 
		"0000000111000000", 
		"0000000111000000", 
		"0000000111000000", 
		"0000000111000000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_score_2	: array_16x16 :=
		("0000000000000000", --2 used for keeping score
		"0000000000000000", 
		"0000000000000000", 
		"0000111111110000", 
		"0001111111111000", 
		"0001110000111000", 
		"0000000000111000", 
		"0000000001110000", 
		"0000000011100000", 
		"0000000111000000", 
		"0000001110000000", 
		"0000111111111000", 
		"0001111111111000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_score_3	: array_16x16 :=
		("0000000000000000", --3 used for keeping score
		"0000000000000000", 
		"0000000000000000", 
		"0000111111110000", 
		"0001111111111000", 
		"0001100000011000", 
		"0000000000011000", 
		"0000000111110000", 
		"0000000111110000", 
		"0000000000011000", 
		"0001100000011000", 
		"0001111111111000", 
		"0000111111110000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_score_4	: array_16x16 :=
		("0000000000000000", --4 used for keepig score
		"0000000000000000", 
		"0000000000000000", 
		"0000000011111000", 
		"0000000111111000", 
		"0000001110011000", 
		"0000011100011000", 
		"0000111000011000", 
		"0001111111111100", 
		"0001111111111100", 
		"0000000000011000", 
		"0000000000011000", 
		"0000000000011000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_score_5	: array_16x16 :=
		("0000000000000000", --5 used for keeping score
		"0000000000000000", 
		"0000000000000000", 
		"0001111111111000", 
		"0001111111111000", 
		"0001100000000000", 
		"0001100000000000", 
		"0001111111110000", 
		"0001111111111000", 
		"0000000000011000", 
		"0001100000011000", 
		"0001111111111000", 
		"0000111111110000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_score_6	: array_16x16 :=
		("0000000000000000", --6 used for keeping score
		"0000000000000000", 
		"0000000000000000", 
		"0000111111110000", 
		"0001111111111000", 
		"0001100000011000", 
		"0001100000000000", 
		"0001111111110000", 
		"0001111111111000", 
		"0001100000011000", 
		"0001100000011000", 
		"0001111111111000", 
		"0000111111110000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_score_7	: array_16x16 :=
		("0000000000000000", --7 used for keeping score
		"0000000000000000", 
		"0000000000000000", 
		"0001111111111000", 
		"0001111111111000", 
		"0000000001110000", 
		"0000000001110000", 
		"0000000011100000", 
		"0000000011100000", 
		"0000000111000000", 
		"0000000111000000", 
		"0000001110000000", 
		"0000001110000000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_score_8	: array_16x16 :=
		("0000000000000000", --8 used for keeping score
		"0000000000000000", 
		"0000000000000000", 
		"0000111111110000", 
		"0001111111111000", 
		"0001100000011000", 
		"0001100000011000", 
		"0000111111110000", 
		"0000111111110000", 
		"0001100000011000", 
		"0001100000011000", 
		"0001111111111000", 
		"0000111111110000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	constant sprite_score_9	: array_16x16 :=
		("0000000000000000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000111111110000", 
		"0001111111111000", 
		"0001100000011000", 
		"0001100000011000", 
		"0001111111111000", 
		"0000111111111000", 
		"0000000000011000", 
		"0001100000011000", 
		"0001111111111000", 
		"0000111111110000", 
		"0000000000000000", 
		"0000000000000000", 
		"0000000000000000");
	
	
	signal sprite_2 : img;
	signal sprite_4 : img;
	signal sprite_8 : img;
	signal sprite_16 : img;
	signal sprite_32 : img;
	signal sprite_64 : img;
	signal sprite_128 : img;
	signal sprite_256 : img;
	signal sprite_512 : img;
	signal sprite_1024 : img;
	signal sprite_2048 : img;
	
	
	--signal sprite_sel : std_logic_vector (3 downto 0) := "0001";--take out later, just for testing 2
	
	Begin
		
		
		--in game
		--sprites yo
		--booyah
		--reminder to make another process for sending out the other sprites
		--leave the top 6 blank and bottom 6 blank
		
		
		sprite_2(0)			<="000000000000000000000000000000000000000000000000";
		sprite_2(1)			<="000000000000000000000000000000000000000000000000";
		sprite_2(2)			<="000000000000000000000000000000000000000000000000";
		sprite_2(3)			<="000000000000000000000000000000000000000000000000";
		sprite_2(4)			<="000000000000000000000000000000000000000000000000";
		sprite_2(5)			<="000000000000000001111111111111111000000000000000";
		sprite_2(6)			<="000000000000001111111111111111111111000000000000";
		sprite_2(7)			<="000000000000011111111111111111111111100000000000";
		sprite_2(8)			<="000000000000011111110000000000111111100000000000";
		sprite_2(9)			<="000000000000000000000000000001111111000000000000";
		sprite_2(10)		<="000000000000000000000000000011111110000000000000";
		sprite_2(11)		<="000000000000000000000000000111111100000000000000";
		sprite_2(12)		<="000000000000000000000000001111111000000000000000";
		sprite_2(13)		<="000000000000000000000000011111110000000000000000";
		sprite_2(14)		<="000000000000000000000000111111100000000000000000";
		sprite_2(15)		<="000000000000000000000001111111000000000000000000";
		sprite_2(16)		<="000000000000000000000011111110000000000000000000";
		sprite_2(17)		<="000000000000000000000111111100000000000000000000";
		sprite_2(18)		<="000000000000000000001111111000000000000000000000";
		sprite_2(19)		<="000000000000000000011111110000000000000000000000";
		sprite_2(20)		<="000000000000000000111111100000000000000000000000";
		sprite_2(21)		<="000000000000000001111111000000000000000000000000";
		sprite_2(22)		<="000000000000000011111111000000000000000000000000";
		sprite_2(23)		<="000000000000001111111110000000000000000000000000";
		sprite_2(24)		<="000000000000111111111111111111111111100000000000";
		sprite_2(25)		<="000000000000111111111111111111111111100000000000";
		sprite_2(26)		<="000000000000000000000000000000000000000000000000";
		sprite_2(27)		<="000000000000000000000000000000000000000000000000";
		sprite_2(28)		<="000000000000000000000000000000000000000000000000";
		sprite_2(29)		<="000000000000000000000000000000000000000000000000";
		sprite_2(30)		<="000000000000000000000000000000000000000000000000";
		sprite_2(31)		<="000000000000000000000000000000000000000000000000";
		
		
		
		sprite_4(0)			<="000000000000000000000000000000000000000000000000";
		sprite_4(1)			<="000000000000000000000000000000000000000000000000";
		sprite_4(2)			<="000000000000000000000000000000000000000000000000";
		sprite_4(3)			<="000000000000000000000000000000000000000000000000";
		sprite_4(4)			<="000000000000000000000000000000000000000000000000";
		sprite_4(5)			<="000000000000000000000000000000000000000000000000";
		sprite_4(6)			<="000000000000000000000000111111111111000000000000";
		sprite_4(7)			<="000000000000000000000001111111111111000000000000";
		sprite_4(8)			<="000000000000000000000011111100011111000000000000";
		sprite_4(9)			<="000000000000000000000111111000011111000000000000";
		sprite_4(10)		<="000000000000000000001111110000011111000000000000";
		sprite_4(11)		<="000000000000000000011111100000011111000000000000";
		sprite_4(12)		<="000000000000000000111111000000011111000000000000";
		sprite_4(13)		<="000000000000000001111110000000011111000000000000";
		sprite_4(14)		<="000000000000000011111100000000011111000000000000";
		sprite_4(15)		<="000000000000000111111000000000011111000000000000";
		sprite_4(16)		<="000000000000001111110000000000011111000000000000";
		sprite_4(17)		<="000000000000011111100000000000011111000000000000";
		sprite_4(18)		<="000000000000111111000000000000011111000000000000";
		sprite_4(19)		<="000000000001111110000000000000011111000000000000";
		sprite_4(20)		<="000000000011111111111111111111111111110000000000";
		sprite_4(21)		<="000000000111111111111111111111111111110000000000";
		sprite_4(22)		<="000000000011111111111111111111111111100000000000";
		sprite_4(23)		<="000000000000000000000000000000011111000000000000";
		sprite_4(24)		<="000000000000000000000000000000011111000000000000";
		sprite_4(25)		<="000000000000000000000000000000011111000000000000";
		sprite_4(26)		<="000000000000000000000000000000011111000000000000";
		sprite_4(27)		<="000000000000000000000000000000000000000000000000";
		sprite_4(28)		<="000000000000000000000000000000000000000000000000";
		sprite_4(29)		<="000000000000000000000000000000000000000000000000";
		sprite_4(30)		<="000000000000000000000000000000000000000000000000";
		sprite_4(31)		<="000000000000000000000000000000000000000000000000";
		
		
		
		sprite_8(0)			<="000000000000000000000000000000000000000000000000";
		sprite_8(1)			<="000000000000000000000000000000000000000000000000";
		sprite_8(2)			<="000000000000000000000000000000000000000000000000";
		sprite_8(3)			<="000000000000000000000000000000000000000000000000";
		sprite_8(4)			<="000000000000000000001111111111000000000000000000";
		sprite_8(5)			<="000000000000000001111111111111111000000000000000";
		sprite_8(6)			<="000000000000001111111111111111111111000000000000";
		sprite_8(7)			<="000000000000011111111100000011111111100000000000";
		sprite_8(8)			<="000000000000111111110000000000111111110000000000";
		sprite_8(9)			<="000000000000111111100000000000011111110000000000";
		sprite_8(10)		<="000000000000111111100000000000011111110000000000";
		sprite_8(11)		<="000000000000111111110000000000111111110000000000";
		sprite_8(12)		<="000000000000011111110000000000111111100000000000";
		sprite_8(13)		<="000000000000001111111000000001111111000000000000";
		sprite_8(14)		<="000000000000000111111111111111111110000000000000";
		sprite_8(15)		<="000000000000000011111111111111111100000000000000";
		sprite_8(16)		<="000000000000000111111111111111111110000000000000";
		sprite_8(17)		<="000000000000001111111000000001111111000000000000";
		sprite_8(18)		<="000000000000011111111000000001111111100000000000";
		sprite_8(19)		<="000000000000111111110000000000111111110000000000";
		sprite_8(20)		<="000000000000111111100000000000011111110000000000";
		sprite_8(21)		<="000000000000111111100000000000011111110000000000";
		sprite_8(22)		<="000000000000011111100000000000011111100000000000";
		sprite_8(23)		<="000000000000011111111000000001111111100000000000";
		sprite_8(24)		<="000000000000001111111111111111111111000000000000";
		sprite_8(25)		<="000000000000000001111111111111111100000000000000";
		sprite_8(26)		<="000000000000000000001111111111110000000000000000";
		sprite_8(27)		<="000000000000000000000000000000000000000000000000";
		sprite_8(28)		<="000000000000000000000000000000000000000000000000";
		sprite_8(29)		<="000000000000000000000000000000000000000000000000";
		sprite_8(30)		<="000000000000000000000000000000000000000000000000";
		sprite_8(31)		<="000000000000000000000000000000000000000000000000";
		
		
		sprite_16(0)			<="000000000000000000000000000000000000000000000000";
		sprite_16(1)			<="000000000000000000000000000000000000000000000000";
		sprite_16(2)			<="000000000000000000000000000000000000000000000000";
		sprite_16(3)			<="000000000000000000000000000000000000000000000000";
		sprite_16(4)			<="000000000000000000000000000000000000000000000000";
		sprite_16(5)			<="000000000000000000000000000000000000000000000000";
		sprite_16(6)			<="000000011111000000000000000000000001111100000000";
		sprite_16(7)			<="000000111111000000000000000000000111111000000000";
		sprite_16(8)			<="000001111111000000000000000000001111110000000000";
		sprite_16(9)			<="000011111111000000000000000000011111100000000000";
		sprite_16(10)			<="000111111111000000000000000000111111000000000000";
		sprite_16(11)			<="000000011111000000000000000001111110000000000000";
		sprite_16(12)			<="000000011111000000000000000011111100000000000000";
		sprite_16(13)			<="000000011111000000000000000111111000000000000000";
		sprite_16(14)			<="000000011111000000000000011111110000000000000000";
		sprite_16(15)			<="000000011111000000000001111111100000000000000000";
		sprite_16(16)			<="000000011111000000000011111111000000000000000000";
		sprite_16(17)			<="000000011111000000001111111111111110000000000000";
		sprite_16(18)			<="000000011111000000011111110000011111110000000000";
		sprite_16(19)			<="000000011111000000111111000000000111111000000000";
		sprite_16(20)			<="000000011111000001111111000000000111111100000000";
		sprite_16(21)			<="000000011111000011111110000000000011111110000000";
		sprite_16(22)			<="000000011111000011111111000000000111111110000000";
		sprite_16(23)			<="000000011111000001111111100000001111111100000000";
		sprite_16(24)			<="000000011111000000111111111111111111111000000000";
		sprite_16(25)			<="000000011111000000001111111111111111110000000000";
		sprite_16(26)			<="000000011111000000000001111111111111000000000000";
		sprite_16(27)			<="000000000000000000000000000000000000000000000000";
		sprite_16(28)			<="000000000000000000000000000000000000000000000000";
		sprite_16(29)			<="000000000000000000000000000000000000000000000000";
		sprite_16(30)			<="000000000000000000000000000000000000000000000000";
		sprite_16(31)			<="000000000000000000000000000000000000000000000000";
		
		
		sprite_32(0)			<="000000000000000000000000000000000000000000000000";
		sprite_32(1)			<="000000000000000000000000000000000000000000000000";
		sprite_32(2)			<="000000000000000000000000000000000000000000000000";
		sprite_32(3)			<="000000000000000000000000000000000000000000000000";
		sprite_32(4)			<="000000000000000000000000000000000000000000000000";
		sprite_32(5)			<="000000000000000000000000000000000000000000000000";
		sprite_32(6)			<="000000111111111111100000000000001111111111100000";
		sprite_32(7)			<="000011111111111111111100000000111111111111111100";
		sprite_32(8)			<="000111111000000001111110000001111110000001111100";
		sprite_32(9)			<="001111100000000001111111000011111000000001111100";
		sprite_32(10)			<="000000000000000001111111000000000000000011111000";
		sprite_32(11)			<="000000000000000011111110000000000000000111111000";
		sprite_32(12)			<="000000000000000111111110000000000000001111110000";
		sprite_32(13)			<="000000000000001111111100000000000000011111100000";
		sprite_32(14)			<="000000001111111111111100000000000000111111000000";
		sprite_32(15)			<="000000001111111111111000000000000001111110000000";
		sprite_32(16)			<="000000001111111111111100000000000011111100000000";
		sprite_32(17)			<="000000000000000111111110000000000111111000000000";
		sprite_32(18)			<="000000000000000011111110000000001111110000000000";
		sprite_32(19)			<="000000000000000001111111000000011111100000000000";
		sprite_32(20)			<="000000000000000000111111000000111111000000000000";
		sprite_32(21)			<="000000000000000001111111000001111110000000000000";
		sprite_32(22)			<="000000000000000011111110000011111100000000000000";
		sprite_32(23)			<="000111110000000111111100000111111110000000000000";
		sprite_32(24)			<="000011111111111111111000000111111111111111111100";
		sprite_32(25)			<="000000111111111111110000000111111111111111111100";
		sprite_32(26)			<="000000000000000000000000000000000000000000000000";
		sprite_32(27)			<="000000000000000000000000000000000000000000000000";
		sprite_32(28)			<="000000000000000000000000000000000000000000000000";
		sprite_32(29)			<="000000000000000000000000000000000000000000000000";
		sprite_32(30)			<="000000000000000000000000000000000000000000000000";
		sprite_32(31)			<="000000000000000000000000000000000000000000000000";

		
		
		sprite_64(0)			<="000000000000000000000000000000000000000000000000";
		sprite_64(1)			<="000000000000000000000000000000000000000000000000";
		sprite_64(2)			<="000000000000000000000000000000000000000000000000";
		sprite_64(3)			<="000000000000000000000000000000000000000000000000";
		sprite_64(4)			<="000000000000000000000000000000000000000000000000";
		sprite_64(5)			<="000000000000000000000000000000000000000000000000";
		sprite_64(6)			<="000000000000000011111000000000000000111111110000";
		sprite_64(7)			<="000000000000000111110000000000000001111111110000";
		sprite_64(8)			<="000000000000001111100000000000000111111111110000";
		sprite_64(9)			<="000000000000111111000000000000000111100111110000";
		sprite_64(10)			<="000000000001111100000000000000001111000111110000";
		sprite_64(11)			<="000000000011111000000000000000011110000111110000";
		sprite_64(12)			<="000000000111111000000000000000111100000111110000";
		sprite_64(13)			<="000000001111110000000000000000111100000111110000";
		sprite_64(14)			<="000000011111100000000000000001111000000111110000";
		sprite_64(15)			<="000001111111000000000000000011111000000111110000";
		sprite_64(16)			<="000011111110000000000000000111110000000111110000";
		sprite_64(17)			<="000011111111111111000000000111110000000111110000";
		sprite_64(18)			<="000111110000001111110000001111100000000111110000";
		sprite_64(19)			<="001111110000000111111000011111111111111111111100";
		sprite_64(20)			<="011111100000000011111100011111111111111111111100";
		sprite_64(21)			<="011111100000000011111100000000000000000111110000";
		sprite_64(22)			<="001111110000000111111000000000000000000111110000";
		sprite_64(23)			<="000111111000000111111000000000000000000111110000";
		sprite_64(24)			<="000011111111111111110000000000000000000111110000";
		sprite_64(25)			<="000000011111111111000000000000000000000111110000";
		sprite_64(26)			<="000000000000000000000000000000000000000000000000";
		sprite_64(27)			<="000000000000000000000000000000000000000000000000";
		sprite_64(28)			<="000000000000000000000000000000000000000000000000";
		sprite_64(29)			<="000000000000000000000000000000000000000000000000";
		sprite_64(30)			<="000000000000000000000000000000000000000000000000";
		sprite_64(31)			<="000000000000000000000000000000000000000000000000";
		
		
		sprite_128(0)			<="000000000000000000000000000000000000000000000000";
		sprite_128(1)			<="000000000000000000000000000000000000000000000000";
		sprite_128(2)			<="000000000000000000000000000000000000000000000000";
		sprite_128(3)			<="000000000000000000000000000000000000000000000000";
		sprite_128(4)			<="000000000000000000000000000000000000000000000000";
		sprite_128(5)			<="000000000000000000000000000000000000000000000000";
		sprite_128(6)			<="000000000000000000000000000000000000000000000000";
		sprite_128(7)			<="000000000000000000000000000000000000000000000000";
		sprite_128(8)			<="000000000000000000111111100000000011111111110000";
		sprite_128(9)			<="000011111000000111111111111000001111111111111000";
		sprite_128(10)			<="000111111000011110000000111100011111100001111100";
		sprite_128(11)			<="001111111000111100000000111100011111000000111100";
		sprite_128(12)			<="000000111000000000000001111000011111000000111100";
		sprite_128(13)			<="000000111000000000000011110000001111100001111000";
		sprite_128(14)			<="000000111000000000000111100000000111111111110000";
		sprite_128(15)			<="000000111000000000001111000000000111111111110000";
		sprite_128(16)			<="000000111000000000011110000000001111100001111000";
		sprite_128(17)			<="000000111000000000111100000000011111000000111100";
		sprite_128(18)			<="000000111000000001111000000000111110000000111110";
		sprite_128(19)			<="000000111000000011110000000000111110000000111110";
		sprite_128(20)			<="000000111000000111100000000000011111000000111100";
		sprite_128(21)			<="000000111000001111000000000000001111100001111000";
		sprite_128(22)			<="000000111000011111111111111111000111111111110000";
		sprite_128(23)			<="000000111000011111111111111111000001111111100000";
		sprite_128(24)			<="000000000000000000000000000000000000000000000000";
		sprite_128(25)			<="000000000000000000000000000000000000000000000000";
		sprite_128(26)			<="000000000000000000000000000000000000000000000000";
		sprite_128(27)			<="000000000000000000000000000000000000000000000000";
		sprite_128(28)			<="000000000000000000000000000000000000000000000000";
		sprite_128(29)			<="000000000000000000000000000000000000000000000000";
		sprite_128(30)			<="000000000000000000000000000000000000000000000000";
		sprite_128(31)			<="000000000000000000000000000000000000000000000000";

		
		
		sprite_256(0)			<="000000000000000000000000000000000000000000000000";
		sprite_256(1)			<="000000000000000000000000000000000000000000000000";
		sprite_256(2)			<="000000000000000000000000000000000000000000000000";
		sprite_256(3)			<="000000000000000000000000000000000000000000000000";
		sprite_256(4)			<="000000000000000000000000000000000000000000000000";
		sprite_256(5)			<="000000000000000000000000000000000000000000000000";
		sprite_256(6)			<="000000000000000000000000000000000000000000000000";
		sprite_256(7)			<="000000000000000000000000000000000000000000000000";
		sprite_256(8)			<="000000111111111000011111111111100000000000111100";
		sprite_256(9)			<="000011111111111110011111111111100000000001111000";
		sprite_256(10)			<="000111100000011110011110000000000000000011110000";
		sprite_256(11)			<="011110000000111100011110000000000000000111100000";
		sprite_256(12)			<="000000000001111000011110000000000000001111000000";
		sprite_256(13)			<="000000000011110000011110000000000000011110000000";
		sprite_256(14)			<="000000000111100000011110000000000000111100000000";
		sprite_256(15)			<="000000001111000000000111111100000001111000000000";
		sprite_256(16)			<="000000011110000000000000011111000011111111000000";
		sprite_256(17)			<="000000111100000000000000000011110111110111110000";
		sprite_256(18)			<="000001111000000000000000000011110111100001111000";
		sprite_256(19)			<="000011110000000000000000000111100111100000111100";
		sprite_256(20)			<="000111100000000000000000001111000111100000111100";
		sprite_256(21)			<="001111111111111100000000111111000011110001111000";
		sprite_256(22)			<="001111111111111100011111111000000000111111100000";
		sprite_256(23)			<="000000000000000000000000000000000000000000000000";
		sprite_256(24)			<="000000000000000000000000000000000000000000000000";
		sprite_256(25)			<="000000000000000000000000000000000000000000000000";
		sprite_256(26)			<="000000000000000000000000000000000000000000000000";
		sprite_256(27)			<="000000000000000000000000000000000000000000000000";
		sprite_256(28)			<="000000000000000000000000000000000000000000000000";
		sprite_256(29)			<="000000000000000000000000000000000000000000000000";
		sprite_256(30)			<="000000000000000000000000000000000000000000000000";
		sprite_256(31)			<="000000000000000000000000000000000000000000000000";
		
		
		
		sprite_512(0)			<="000000000000000000000000000000000000000000000000";
		sprite_512(1)			<="000000000000000000000000000000000000000000000000";
		sprite_512(2)			<="000000000000000000000000000000000000000000000000";
		sprite_512(3)			<="000000000000000000000000000000000000000000000000";
		sprite_512(4)			<="000000000000000000000000000000000000000000000000";
		sprite_512(5)			<="000000000000000000000000000000000000000000000000";
		sprite_512(6)			<="000000000000000000000000000000000000000000000000";
		sprite_512(7)			<="000000000000000000000000000000000001111111100000";
		sprite_512(8)			<="000001111111111110000011110000000111111111111000";
		sprite_512(9)			<="000011111111111110001111110000011110000000111100";
		sprite_512(10)			<="000011110000000000011111110000111100000000111100";
		sprite_512(11)			<="000011110000000000000011110000000000000001111000";
		sprite_512(12)			<="000011110000000000000011110000000000000011110000";
		sprite_512(13)			<="000011110000000000000011110000000000000111100000";
		sprite_512(14)			<="000011110000000000000011110000000000001111000000";
		sprite_512(15)			<="000000111110000000000011110000000000011110000000";
		sprite_512(16)			<="000000000111110000000011110000000000111100000000";
		sprite_512(17)			<="000000000001111100000011110000000001111000000000";
		sprite_512(18)			<="000000000000111110000011110000000011110000000000";
		sprite_512(19)			<="000000000000111100000011110000000111100000000000";
		sprite_512(20)			<="000000000011110000000011110000001111111111111000";
		sprite_512(21)			<="000011111111100000000011110000001111111111111000";
		sprite_512(22)			<="000000000000000000000000000000000000000000000000";
		sprite_512(23)			<="000000000000000000000000000000000000000000000000";
		sprite_512(24)			<="000000000000000000000000000000000000000000000000";
		sprite_512(25)			<="000000000000000000000000000000000000000000000000";
		sprite_512(26)			<="000000000000000000000000000000000000000000000000";
		sprite_512(27)			<="000000000000000000000000000000000000000000000000";
		sprite_512(28)			<="000000000000000000000000000000000000000000000000";
		sprite_512(29)			<="000000000000000000000000000000000000000000000000";
		sprite_512(30)			<="000000000000000000000000000000000000000000000000";
		sprite_512(31)			<="000000000000000000000000000000000000000000000000";

		
		
		sprite_1024(0)			<="000000000000000000000000000000000000000000000000";
		sprite_1024(1)			<="000000000000000000000000000000000000000000000000";
		sprite_1024(2)			<="000000000000111100000000000000111110000000000000";
		sprite_1024(3)			<="000000000011111100000000000011111111100000000000";
		sprite_1024(4)			<="000000000111111100000000001111111111111000000000";
		sprite_1024(5)			<="000000001111111100000000011111000000111100000000";
		sprite_1024(6)			<="000000000000111100000000111110000000011110000000";
		sprite_1024(7)			<="000000000000111100000000111100000000011110000000";
		sprite_1024(8)			<="000000000000111100000000111100000000011110000000";
		sprite_1024(9)			<="000000000000111100000000111100000000011110000000";
		sprite_1024(10)		<="000000000000111100000000111100000000011110000000";
		sprite_1024(11)		<="000000000000111100000000111100000000011110000000";
		sprite_1024(12)		<="000000000000111100000000011111000000111100000000";
		sprite_1024(13)		<="000000000000111100000000001111111111111000000000";
		sprite_1024(14)		<="000000000000111100000000000001111111100000000000";
		sprite_1024(15)		<="000000000000000000000000000000000000000000000000";
		sprite_1024(16)		<="000000000011111111100000000000001111110000000000";
		sprite_1024(17)		<="000000001111111111111000000000011111110000000000";
		sprite_1024(18)		<="000000011110000001111000000000111111110000000000";
		sprite_1024(19)		<="000000000000000001111000000011110011110000000000";
		sprite_1024(20)		<="000000000000000011110000000111100011110000000000";
		sprite_1024(21)		<="000000000000000111100000001111000011110000000000";
		sprite_1024(22)		<="000000000000001111000000011110000011110000000000";
		sprite_1024(23)		<="000000000000011110000000111100000011110000000000";
		sprite_1024(24)		<="000000000000111100000001111000000011110000000000";
		sprite_1024(25)		<="000000000001111000000011111111111111111000000000";
		sprite_1024(26)		<="000000000011110000000011111111111111111000000000";
		sprite_1024(27)		<="000000000111100000000000000000000011110000000000";
		sprite_1024(28)		<="000000001111111111111000000000000011110000000000";
		sprite_1024(29)		<="000000001111111111111000000000000011110000000000";
		sprite_1024(30)		<="000000000000000000000000000000000000000000000000";
		sprite_1024(31)		<="000000000000000000000000000000000000000000000000";
		
		
		sprite_2048(0)			<="000000000000000000000000000000000000000000000000";
		sprite_2048(1)			<="000000011111111111000000000001111111111100000000";
		sprite_2048(2)			<="000001111111111111100000000111111000111110000000";
		sprite_2048(3)			<="000011110000000111100000001111000000001111000000";
		sprite_2048(4)			<="000000000000000111100000011111000000001111100000";
		sprite_2048(5)			<="000000000000001111000000011111000000001111100000";
		sprite_2048(6)			<="000000000000011110000000011110000000000111100000";
		sprite_2048(7)			<="000000000000111100000000011110000000000111100000";
		sprite_2048(8)			<="000000000001111000000000011110000000000111100000";
		sprite_2048(9)			<="000000000011110000000000011110000000000111100000";
		sprite_2048(10)		<="000000000111100000000000011111000000001111100000";
		sprite_2048(11)		<="000000001111000000000000001111000000001111000000";
		sprite_2048(12)		<="000000011110000000000000001111000000001111000000";
		sprite_2048(13)		<="000000111100000000000000000111111000111110000000";
		sprite_2048(14)		<="000001111111111111000000000001111111111000000000";
		sprite_2048(15)		<="000001111111111111000000000000011111100000000000";
		sprite_2048(16)		<="000000000000000000000000000000000000000000000000";
		sprite_2048(17)		<="000000000001111110000000000000011111110000000000";
		sprite_2048(18)		<="000000000011111110000000000001111111111100000000";
		sprite_2048(19)		<="000000000111111110000000000011110000011110000000";
		sprite_2048(20)		<="000000011110011110000000000011110000011110000000";
		sprite_2048(21)		<="000000111100011110000000000001111000111100000000";
		sprite_2048(22)		<="000001111000011110000000000001111111111100000000";
		sprite_2048(23)		<="000011110000011110000000000001111111111100000000";
		sprite_2048(24)		<="000111100000011110000000000011110000011110000000";
		sprite_2048(25)		<="001111000000011110000000000111100000001111000000";
		sprite_2048(26)		<="011111111111111111000000000111100000001111000000";
		sprite_2048(27)		<="011111111111111111000000000011110000011110000000";
		sprite_2048(28)		<="000000000000011110000000000001111000111100000000";
		sprite_2048(29)		<="000000000000011110000000000000011111111000000000";
		sprite_2048(30)		<="000000000000011110000000000000000111100000000000";
		sprite_2048(31)		<="000000000000000000000000000000000000000000000000";


		
		
		
		Sprite_out_score : process(DrawX, DrawY, scoreIn)
		begin
			--DrawX >= 520 and DrawX <= 620 and DrawY >= 220 and DrawY <= 260
			if (DrawX >= 525 and DrawX <= 540 and DrawY >= 222 and DrawY <= 237) then
				score_sprite_out <= sprite_S;
			elsif (DrawX >= 542 and DrawX <= 557 and DrawY >= 222 and DrawY <= 237) then
				score_sprite_out <= sprite_C;
			elsif (DrawX >= 559 and DrawX <= 574 and DrawY >= 222 and DrawY <= 237) then
				score_sprite_out <= sprite_O;
			elsif (DrawX >= 576 and DrawX <= 591 and DrawY >= 222 and DrawY <= 237) then
				score_sprite_out <= sprite_R;
			elsif (DrawX >= 593 and DrawX <= 608 and DrawY >= 222 and DrawY <= 237) then
				score_sprite_out <= sprite_E;
			--now for score numbers
			elsif (DrawX >= 525 and DrawX <= 540 and DrawY >= 240 and DrawY <= 255) then
				if (scoreIn(4) = 0) then
					score_sprite_out <= sprite_score_0;
				elsif (scoreIn(4) = 1) then
					score_sprite_out <= sprite_score_1;
				elsif (scoreIn(4) = 2) then
					score_sprite_out <= sprite_score_2;
				elsif (scoreIn(4) = 3) then
					score_sprite_out <= sprite_score_3;
				elsif (scoreIn(4) = 4) then
					score_sprite_out <= sprite_score_4;
				elsif (scoreIn(4) = 5) then
					score_sprite_out <= sprite_score_5;
				elsif (scoreIn(4) = 6) then
					score_sprite_out <= sprite_score_6;
				elsif (scoreIn(4) = 7) then
					score_sprite_out <= sprite_score_7;
				elsif (scoreIn(4) = 8) then
					score_sprite_out <= sprite_score_8;
				elsif (scoreIn(4) = 9) then
					score_sprite_out <= sprite_score_9;
				else
					score_sprite_out <= sprite_score_0;
				end if;
			elsif (DrawX >= 542 and DrawX <= 557 and DrawY >= 240 and DrawY <= 255) then
				if (scoreIn(3) = 0) then
					score_sprite_out <= sprite_score_0;
				elsif (scoreIn(3) = 1) then
					score_sprite_out <= sprite_score_1;
				elsif (scoreIn(3) = 2) then
					score_sprite_out <= sprite_score_2;
				elsif (scoreIn(3) = 3) then
					score_sprite_out <= sprite_score_3;
				elsif (scoreIn(3) = 4) then
					score_sprite_out <= sprite_score_4;
				elsif (scoreIn(3) = 5) then
					score_sprite_out <= sprite_score_5;
				elsif (scoreIn(3) = 6) then
					score_sprite_out <= sprite_score_6;
				elsif (scoreIn(3) = 7) then
					score_sprite_out <= sprite_score_7;
				elsif (scoreIn(3) = 8) then
					score_sprite_out <= sprite_score_8;
				elsif (scoreIn(3) = 9) then
					score_sprite_out <= sprite_score_9;
				else
					score_sprite_out <= sprite_score_0;
				end if;
			elsif (DrawX >= 559 and DrawX <= 574 and DrawY >= 240 and DrawY <= 255) then
				if (scoreIn(2) = 0) then
					score_sprite_out <= sprite_score_0;
				elsif (scoreIn(2) = 1) then
					score_sprite_out <= sprite_score_1;
				elsif (scoreIn(2) = 2) then
					score_sprite_out <= sprite_score_2;
				elsif (scoreIn(2) = 3) then
					score_sprite_out <= sprite_score_3;
				elsif (scoreIn(2) = 4) then
					score_sprite_out <= sprite_score_4;
				elsif (scoreIn(2) = 5) then
					score_sprite_out <= sprite_score_5;
				elsif (scoreIn(2) = 6) then
					score_sprite_out <= sprite_score_6;
				elsif (scoreIn(2) = 7) then
					score_sprite_out <= sprite_score_7;
				elsif (scoreIn(2) = 8) then
					score_sprite_out <= sprite_score_8;
				elsif (scoreIn(2) = 9) then
					score_sprite_out <= sprite_score_9;
				else
					score_sprite_out <= sprite_score_0;
				end if;
			elsif (DrawX >= 576 and DrawX <= 591 and DrawY >= 240 and DrawY <= 255) then
				if (scoreIn(1) = 0) then
					score_sprite_out <= sprite_score_0;
				elsif (scoreIn(1) = 1) then
					score_sprite_out <= sprite_score_1;
				elsif (scoreIn(1) = 2) then
					score_sprite_out <= sprite_score_2;
				elsif (scoreIn(1) = 3) then
					score_sprite_out <= sprite_score_3;
				elsif (scoreIn(1) = 4) then
					score_sprite_out <= sprite_score_4;
				elsif (scoreIn(1) = 5) then
					score_sprite_out <= sprite_score_5;
				elsif (scoreIn(1) = 6) then
					score_sprite_out <= sprite_score_6;
				elsif (scoreIn(1) = 7) then
					score_sprite_out <= sprite_score_7;
				elsif (scoreIn(1) = 8) then
					score_sprite_out <= sprite_score_8;
				elsif (scoreIn(1) = 9) then
					score_sprite_out <= sprite_score_9;
				else
					score_sprite_out <= sprite_score_3;
				end if;
			elsif (DrawX >= 593 and DrawX <= 608 and DrawY >= 240 and DrawY <= 255) then
				if (scoreIn(0) = 0) then
					score_sprite_out <= sprite_score_0;
				elsif (scoreIn(0) = 1) then
					score_sprite_out <= sprite_score_1;
				elsif (scoreIn(0) = 2) then
					score_sprite_out <= sprite_score_2;
				elsif (scoreIn(0) = 3) then
					score_sprite_out <= sprite_score_3;
				elsif (scoreIn(0) = 4) then
					score_sprite_out <= sprite_score_4;
				elsif (scoreIn(0) = 5) then
					score_sprite_out <= sprite_score_5;
				elsif (scoreIn(0) = 6) then
					score_sprite_out <= sprite_score_6;
				elsif (scoreIn(0) = 7) then
					score_sprite_out <= sprite_score_7;
				elsif (scoreIn(0) = 8) then
					score_sprite_out <= sprite_score_8;
				elsif (scoreIn(0) = 9) then
					score_sprite_out <= sprite_score_9;
				else
					score_sprite_out <= sprite_score_0;
				end if;
			else
				score_sprite_out <= sprite_score_0;
			end if;
			
			
	end process Sprite_out_score;
	--score_sprite_out <= sprite_S;
	--end process;
	
	--sprite_num_color
	--sprite_back_color
	--begin
	sprite_color_intro : process(outSprites, outFree, drawX, drawY, Reset) --trouble getting this to compile -___- lso |||||||||| initial testing run w/2 blocks
		--begin
			variable r : std_logic_vector (9 downto 0) := "0000000000"; --background color
			variable g : std_logic_vector (9 downto 0) := "0000000000";
			variable b : std_logic_vector (9 downto 0) := "0000000000";
			
			variable r_num : std_logic_vector (9 downto 0) := "0000000000"; --number color
			variable g_num : std_logic_vector (9 downto 0) := "0000000000";
			variable b_num : std_logic_vector (9 downto 0) := "0000000000";
			
			variable x : integer range 0 to 3 := 0;
			variable y : integer range 0 to 3 := 0;
			
			begin
			--if (reset = '1') then
					if(DrawX >= 16 and DrawX <= 116 and DrawY >= 16 and DrawY <= 116) then
						x := 0;
						y := 0;
					elsif(DrawX >= 132 and DrawX <= 232 and DrawY >= 16 and DrawY <= 116) then --ifDrawX is in tile zero output sprite in tile 0
						x := 1;
						y := 0;
					elsif (DrawX >= 248 and DrawX <= 348 and DrawY >= 16 and DrawY <= 116) then
						x := 2;
						y := 0;
					elsif (DrawX >= 364 and DrawX <= 464 and DrawY >= 16 and DrawY <= 116) then
						x := 3;
						y := 0;
					elsif (DrawX >= 16 and DrawX <= 116 and DrawY >= 132 and DrawY <= 232) then
						x := 0;
						y := 1;
					elsif (DrawX >= 132 and DrawX <= 232 and DrawY >= 132 and DrawY <= 232) then
						x := 1;
						y := 1;
					elsif (DrawX >= 248 and DrawX <= 348 and DrawY >= 132 and DrawY <= 232) then
						x := 2;
						y := 1;
					elsif (DrawX >= 364 and DrawX <= 464 and DrawY >= 132 and DrawY <= 232) then
						x := 3;
						y := 1;
					elsif (DrawX >= 16 and DrawX <= 116 and DrawY >= 248 and DrawY <= 348) then
						x := 0;
						y := 2;
					elsif (DrawX >= 132 and DrawX <= 232 and DrawY >= 248 and DrawY <= 348) then
						x := 1;
						y := 2;
					elsif (DrawX >= 248 and DrawX <= 348 and DrawY >= 248 and DrawY <= 348) then
						x := 2;
						y := 2;
					elsif (DrawX >= 364 and DrawX <= 464 and DrawY >= 248 and DrawY <= 348) then
						x := 3;
						y := 2;
					elsif (DrawX >= 16 and DrawX <= 116 and DrawY >= 364 and DrawY <= 464) then
						x := 0;
						y := 3;
					elsif (DrawX >= 132 and DrawX <= 232 and DrawY >= 364 and DrawY <= 464) then
						x := 1;
						y := 3;
					elsif (DrawX >= 248 and DrawX <= 348 and DrawY >= 364 and DrawY <= 464) then
						x := 2;
						y := 3;
					elsif (DrawX >= 364 and DrawX <= 464 and DrawY >= 364 and DrawY <= 464) then
						x := 3;
						y := 3;
					else
						x := 0;
						y := 0;
					end if;
					if (outSprites(y,x) = "0001") then --changed from 0001
						r_num := "0000000000";
						g_num := "0000000000";
						b_num := "0000000000";
					
						r := "1111111100";
						g := "1111111100";
						b := "1111111100";
						tile_sprite_out <= sprite_2;

					elsif (outSprites(y,x) = "0010") then --chaned from 0010
						r_num := "0000000000";
						g_num := "0000000000";
						b_num := "0000000000";
					
						r := "1111000000"; --0011111110
						g := "1111000000"; --0011010000
						b := "1111000000"; --0011000000
						tile_sprite_out <= sprite_4;
					
					elsif (outSprites(y,x) = "0011") then --chaned from 0010
						r_num := "1111111111";
						g_num := "1111111111";
						b_num := "1111111111";
					
						r := "1111010000"; --0011111110
						g := "1010010000"; --0011010000
						b := "0110000000"; --0011000000
						tile_sprite_out <= sprite_8;
					
					elsif (outSprites(y,x) = "0100") then --chaned from 0010
						r_num := "1111111111";
						g_num := "1111111111";
						b_num := "1111111111";
					
						r := "1111010000"; --0011111110
						g := "0101001000"; --0011010000
						b := "0011000000"; --0011000000
						tile_sprite_out <= sprite_16;
					
					elsif (outSprites(y,x) = "0101") then --chaned from 0010
						r_num := "1111111111";
						g_num := "1111111111";
						b_num := "1111111111";
					
						r := "1111010000"; --0011111110
						g := "0101001000"; --0011010000
						b := "0011000000"; --0011000000
						tile_sprite_out <= sprite_32;
					
					elsif (outSprites(y,x) = "0110") then --chaned from 0010
						r_num := "1111111111";
						g_num := "1111111111";
						b_num := "1111111111";
					
						r := "1111111111"; --0011111110
						g := "0000000000"; --0011010000
						b := "0000000000"; --0011000000
						tile_sprite_out <= sprite_64;
					
					elsif (outSprites(y,x) = "0111") then --chaned from 0010
						r_num := "1111111111";
						g_num := "1111111111";
						b_num := "1111111111";
					
						r := "0111111111"; --0011111110
						g := "0111111111"; --0011010000
						b := "0000000000"; --0011000000
						tile_sprite_out <= sprite_128;
					
					elsif (outSprites(y,x) = "1000") then --chaned from 0010
						r_num := "1111111111";
						g_num := "1111111111";
						b_num := "1111111111";
					
						r := "1000000000"; --0011111110
						g := "1000000000"; --0011010000
						b := "0000000000"; --0011000000
						tile_sprite_out <= sprite_256;
					
					elsif (outSprites(y,x) = "1001") then --chaned from 0010
						r_num := "1111111111";
						g_num := "1111111111";
						b_num := "1111111111";
					
						r := "1100000000"; --0011111110
						g := "1100000000"; --0011010000
						b := "0000000000"; --0011000000
						tile_sprite_out <= sprite_512;
					
					elsif (outSprites(y,x) = "1010") then --chaned from 0010
						r_num := "1111111111";
						g_num := "1111111111";
						b_num := "1111111111";
					
						r := "1110000000"; --0011111110
						g := "1110000000"; --0011010000
						b := "0000000000"; --0011000000
						tile_sprite_out <= sprite_1024;
					
					elsif (outSprites(y,x) = "1011") then --chaned from 0010
						r_num := "1111111111";
						g_num := "1111111111";
						b_num := "1111111111";
					
						r := "1111111111"; --0011111110
						g := "1111111111"; --0011010000
						b := "0000000000"; --0011000000
						tile_sprite_out <= sprite_2048;
					
					else
						r_num := "0000000000";
						g_num := "0000000000";
						b_num := "0000000000";
					
						r := "0000000000";
						g := "1000000000";
						b := "0000000000";
						tile_sprite_out <= sprite_2;
					end if;
					sprite_back_color <= r & g & b;
					sprite_num_color <= r_num & g_num & b_num;
			--sprite_back_color2 <= r2 & g2 & b2;
			--sprite_num_color2 <= r2_num & g2_num & b2_num;
			--sprite_num_color <= r_num & g_num & b_num;
			--sprite_back_color <= r & g & b;
			--end if;
			--else -- add more for moving
			--end if;
	
	end process sprite_color_intro;
	
	--tile_sprite_out <= sprite_2;




end Behavioral;